`timescale 1ns / 1ps

module mips (
           input clk,
           input reset
       );

endmodule
