

`timescale 1ns / 1ps

module mips (
           input wire clk,
           input wire reset
       );




endmodule
