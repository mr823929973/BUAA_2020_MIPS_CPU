`timescale 1ns / 1ps

module ifu(
           input clk,
           input reset,
           input isBracnch,
           input [31:0] branchAddr,
           input isJump,
           input [31:0] jumpAddr,
           output [31:0] PC,
           output [31:0] instructure
       );



endmodule
