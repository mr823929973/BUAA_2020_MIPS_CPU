`ifndef INSTR_VH
`define INSTR_VH

`define addu 4'd0
`define subu 4'd1
`define ori  4'd2
`define lw   4'd3
`define sw   4'd4
`define beq  4'd5
`define lui  4'd6

`define jal  4'd7
`define jr   4'd8
`define sll  4'd9

`endif